-- ************************************************************************
-- Unified Testbench for ADC (TDC-based and RC-based delta-sigma ADC)
-- Simulates both TDC-based and traditional RC delta-sigma ADC
-- Uses 1.25V effective reference voltage for consistent voltage range, tested empirically in HW
-- ************************************************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library vunit_lib;
context vunit_lib.vunit_context;

library fpga_lib;
use fpga_lib.clk_rst_pkg.all;

entity adc_top_tb is
    generic(
        runner_cfg         : string;
        -- ADC type selection: "tdc" for TDC-based ADC, "rc" for RC delta-sigma ADC
        GC_ADC_TYPE        : string  := "tdc";
        -- Test configuration generics for VUnit
        -- Signal type: 0=sine, 1=DC, 2=ramp, 3=square
        GC_TB_SIGNAL_TYPE  : integer := 0; -- Signal type enum
        GC_TB_AMPLITUDE    : real    := 0.25; -- Signal amplitude (normalized: 0.0 to 1.0, will be scaled to 1.3V)
        GC_TB_FREQUENCY_HZ : real    := 1000.0; -- Frequency for sine/square waves
        GC_TB_DC_LEVEL     : real    := 0.5; -- DC offset or DC test level (normalized: 0.5 = 0.625V at 1.25V reference)
        GC_OPEN_LOOP       : boolean := false -- Enable open-loop mode for DAC characterization
    );
end entity;

architecture behavioral of adc_top_tb is

    -- Test parameters
    constant C_CLK_SYS_PERIOD : time     := 10 ns; -- 100 MHz (from PLL outclk_0 in hardware)
    constant C_CLK_TDC_PERIOD : time     := 2.474 ns; -- 404.166667 MHz (ASYNC from PLL iopll_tdc_outclk0 in hardware)
    constant C_REF_PERIOD     : time     := 20 ns; -- 50 MHz reference (from PLL outclk_2 in hardware)
    constant C_DATA_WIDTH     : positive := 16;
    constant C_TDC_WIDTH      : positive := 16;

    -- DUT signals
    signal clk_sys   : std_logic := '0';
    signal clk_tdc   : std_logic := '0';
    signal reset     : std_logic := '1';
    signal ref_clock : std_logic := '0';

    -- Output signals
    signal sample_data  : std_logic_vector(C_DATA_WIDTH - 1 downto 0);
    signal sample_valid : std_logic;

    -- GPIO IP interface signals
    signal dac_out_bit      : std_logic; -- DAC output from DUT (goes to external RC filter)
    signal s_comparator_out : std_logic_vector(0 downto 0); -- Comparator output (behavioral)

    -- Analog comparator modeling signals
    -- Test realistic power-up conditions: both pins start at same voltage
    -- Initialize to 0V to test worst-case: both inputs equal, no initial differential
    signal analog_voltage_p : real := 0.0; -- P-pin voltage (input signal)
    signal analog_voltage_n : real := 0.0; -- N-pin voltage (from external RC filter)

    -- RC filter internal signals (for ref_clock-rate optimization)
    signal duty_count_reg   : integer range 0 to 255 := 0;
    signal duty_period_done : std_logic              := '0';

    -- Pad-level signals (after threshold conversion)
    signal pad_p : std_logic := '0';    -- P-pad digital (comparator P input)
    signal pad_n : std_logic := '0';    -- N-pad digital (comparator N threshold)

    -- RC ADC comparator signal - simple instantaneous analog comparison
    signal rc_comparator_out : std_logic := '0';

    -- Debug signals for TDC characterization
    signal debug_tdc_out   : signed(C_TDC_WIDTH - 1 downto 0);
    signal debug_tdc_valid : std_logic;
    signal open_loop_dac   : std_logic := '0'; -- Control signal for open-loop tests

    -- Test control
    signal sim_finished    : boolean   := false;
    signal testpoint_reset : std_logic := '0'; -- Pulse to reset TDC monitor between test points
    signal tdc_char_done   : boolean   := false; -- Early termination for TDC characterization

    -- Sample statistics (updated by p_monitor, checked by test process)
    signal sample_min_value : integer := 0;
    signal sample_max_value : integer := 0;
    signal sample_count_sig : integer := 0;
    signal sample_sum_value : integer := 0; -- Sum of all samples for averaging

begin

    -- ========================================================================
    -- Device Under Test - Conditional instantiation based on GC_ADC_TYPE
    -- ========================================================================

    -- TDC ADC instantiation (GC_ADC_TYPE = "tdc")
    g_tdc_adc : if GC_ADC_TYPE = "tdc" generate
        i_dut_tdc : entity work.tdc_adc_top
            generic map(
                GC_DECIMATION => 64,    -- 32us per sample (64 x 500ns) - 6-bit DAC resolution
                GC_DATA_WIDTH => C_DATA_WIDTH,
                GC_TDC_OUTPUT => C_TDC_WIDTH,
                GC_SIM        => false, -- Disable debug reports for fast simulation
                GC_FAST_SIM   => true,  -- Enable fast boot mode (reduced timeouts)
                GC_OPEN_LOOP  => GC_OPEN_LOOP -- Pass through from testbench generic
            )
            port map(
                clk_sys             => clk_sys,
                clk_tdc             => clk_tdc,
                reset               => reset,
                ref_clock           => ref_clock,
                -- GPIO IP interface (real GPIO IP instantiated below)
                comparator_in       => s_comparator_out(0), -- From GPIO IP differential comparator
                dac_out_bit         => dac_out_bit, -- To GPIO DAC IP
                trigger_enable      => '1', -- Always enabled in testbench
                open_loop_dac_duty  => open_loop_dac, -- For characterization tests

                sample_data         => sample_data,
                sample_valid        => sample_valid,
                debug_tdc_out       => debug_tdc_out,
                debug_tdc_valid     => debug_tdc_valid,
                -- TDC monitor outputs (not used in this testbench)
                tdc_monitor_code    => open,
                tdc_monitor_center  => open,
                tdc_monitor_diff    => open,
                tdc_monitor_dac     => open,
                tdc_monitor_valid   => open,
                -- Runtime control (not used in this testbench)
                disable_tdc_contrib => '0',
                disable_eq_filter   => '0',
                disable_lp_filter   => '0'
            );
    end generate;

    -- RC ADC instantiation (GC_ADC_TYPE = "rc")
    g_rc_adc : if GC_ADC_TYPE = "rc" generate
        i_dut_rc : entity work.rc_adc_top
            generic map(
                GC_DECIMATION => 64,    -- Same decimation as TDC for comparison
                GC_DATA_WIDTH => C_DATA_WIDTH
            )
            port map(
                clk          => clk_sys,
                reset        => reset,
                -- Physical ADC interface
                analog_in    => rc_comparator_out, -- From RC-specific comparator model
                dac_out      => dac_out_bit, -- DAC output for feedback
                -- Streaming sample output
                sample_data  => sample_data,
                sample_valid => sample_valid
            );
        -- RC ADC doesn't have TDC debug outputs - tie off
        debug_tdc_out   <= (others => '0');
        debug_tdc_valid <= '0';
    end generate;

    p_behavioral_comparator : process(pad_p, pad_n)
    begin
        -- Differential comparison: pad_p (analog input) vs pad_n (RC filtered feedback)
        -- This matches the actual hardware where comparator compares ANALOG_IN (P-pin)
        -- against ANALOG_IN_N (N-pin, external RC filter from FEEDBACK_OUT)
        if pad_p = '1' and pad_n = '0' then
            s_comparator_out(0) <= '1'; -- Input > Feedback
        elsif pad_p = '0' and pad_n = '1' then
            s_comparator_out(0) <= '0'; -- Input < Feedback
        else
            -- Both same: small signal case, use XOR to create variation
            s_comparator_out(0) <= pad_p xor pad_n;
        end if;
    end process;

    p_clk_sys : process
        variable v_seed1, v_seed2 : positive := 1;
        variable v_rand           : real;
        variable v_init_delay     : time;
    begin
        -- Random initial phase (0 to 5ns) to desynchronize from other clocks
        uniform(v_seed1, v_seed2, v_rand);
        v_init_delay := v_rand * 5.0 ns;
        wait for v_init_delay;

        while not sim_finished loop
            clk_sys <= '0';
            wait for C_CLK_SYS_PERIOD / 2;
            clk_sys <= '1';
            wait for C_CLK_SYS_PERIOD / 2;
        end loop;
        wait;
    end process;

    p_clk_tdc : process
        variable v_seed1, v_seed2 : positive := 2;
        variable v_rand           : real;
        variable v_init_delay     : time;
    begin
        -- Random initial phase (0 to 5ns) to desynchronize from other clocks
        uniform(v_seed1, v_seed2, v_rand);
        v_init_delay := v_rand * 5.0 ns;
        wait for v_init_delay;

        while not sim_finished loop
            clk_tdc <= '0';
            wait for C_CLK_TDC_PERIOD / 2;
            clk_tdc <= '1';
            wait for C_CLK_TDC_PERIOD / 2;
        end loop;
        wait;
    end process;

    p_ref_clock : process
        variable v_seed1, v_seed2 : positive := 3;
        variable v_rand           : real;
        variable v_init_delay     : time;
    begin
        -- Random initial phase (0 to 100ns) to desynchronize from other clocks
        uniform(v_seed1, v_seed2, v_rand);
        v_init_delay := v_rand * 100.0 ns;
        wait for v_init_delay;

        -- Simple reference clock without stress test jitter/ppm
        while not sim_finished loop
            ref_clock <= '0';
            wait for C_REF_PERIOD / 2;

            ref_clock <= '1';
            wait for C_REF_PERIOD / 2;
        end loop;
        wait;
    end process;

    -- ========================================================================
    -- Reset Generation (v8.4: Randomized deassert timing)
    -- ========================================================================
    p_reset : process
        variable v_seed1, v_seed2 : positive := 4;
        variable v_rand           : real;
        variable v_reset_delay    : time;
    begin
        uniform(v_seed1, v_seed2, v_rand);
        v_reset_delay := 200 ns + v_rand * 200 ns;

        reset <= '1';
        wait for v_reset_delay;
        reset <= '0';
        wait;
    end process;

    -- ========================================================================
    -- Analog Signal Generator
    -- ========================================================================
    -- Only update analog value once per ref_clock period instead of every 0.5ns.
    -- This provides massive speedup for AC signals while still being massively
    -- oversampled relative to the 1kHz input frequency.
    -- The comparator/TDC model only samples once per period anyway.
    p_analog_voltage_generator : process
        variable v_time_s : real := 0.0;
        constant C_PI     : real := 3.14159265359;
        constant C_VBANK  : real := 1.25; -- FPGA I/O bank voltage (measured effective Vref)
    begin
        wait until reset = '0';
        report "Analog voltage generator started! Signal type=" & integer'image(GC_TB_SIGNAL_TYPE);

        -- All signal types now update at ref_clock rate (2 MHz)
        -- This is still massively oversampled vs 1kHz input frequency
        loop
            wait until rising_edge(ref_clock);
            v_time_s := v_time_s + real(C_REF_PERIOD / 1 ns) * 1.0e-9;

            case GC_TB_SIGNAL_TYPE is
                when 0 =>               -- Sine wave
                    analog_voltage_p <= (GC_TB_DC_LEVEL + GC_TB_AMPLITUDE * sin(2.0 * C_PI * GC_TB_FREQUENCY_HZ * v_time_s)) * C_VBANK;
                when 1 =>               -- DC level
                    analog_voltage_p <= GC_TB_DC_LEVEL * C_VBANK;
                when 2 =>               -- Ramp (sawtooth)
                    analog_voltage_p <= (GC_TB_DC_LEVEL + GC_TB_AMPLITUDE * (2.0 * ((GC_TB_FREQUENCY_HZ * v_time_s) mod 1.0) - 1.0)) * C_VBANK;
                when 3 =>               -- Square wave
                    if ((GC_TB_FREQUENCY_HZ * v_time_s) mod 1.0) < 0.5 then
                        analog_voltage_p <= (GC_TB_DC_LEVEL + GC_TB_AMPLITUDE) * C_VBANK;
                    else
                        analog_voltage_p <= (GC_TB_DC_LEVEL - GC_TB_AMPLITUDE) * C_VBANK;
                    end if;
                when others =>
                    analog_voltage_p <= 0.0;
            end case;
        end loop;
    end process;

    -- ========================================================================
    -- RC FILTER: Fast ref_clock-rate filter with duty cycle counting
    -- ========================================================================
    -- Duty counter at clk_tdc rate (just counting, no signal updates)
    p_duty_counter : process(clk_tdc, reset)
        constant C_TICKS_PER_PERIOD : integer               := 8; -- 400MHz TDC / 50MHz ref = 8 ticks
        variable v_tick_count       : integer range 0 to 15 := 0;
        variable v_high_count       : integer range 0 to 15 := 0;
    begin
        if reset = '1' then
            v_tick_count     := 0;
            v_high_count     := 0;
            duty_count_reg   <= 0;
            duty_period_done <= '0';
        elsif rising_edge(clk_tdc) then
            -- Count DAC high
            if dac_out_bit = '1' then
                v_high_count := v_high_count + 1;
            end if;
            v_tick_count := v_tick_count + 1;

            -- At end of period, latch count and reset
            if v_tick_count >= C_TICKS_PER_PERIOD then
                duty_count_reg   <= v_high_count;
                duty_period_done <= '1';
                v_tick_count     := 0;
                v_high_count     := 0;
            else
                duty_period_done <= '0';
            end if;
        end if;
    end process;

    -- RC filter at ref_clock rate (only updates when period done)
    p_rc_filter_duty_avg : process(clk_tdc, reset)
        constant C_DAC_HIGH_V       : real      := 1.25;
        constant C_TICKS_PER_PERIOD : integer   := 8; -- 400MHz TDC / 50MHz ref = 8 ticks
        -- RC time constant: tau = 1us (1k x 1nF), T = 20ns (50MHz ref)
        -- alpha = exp(-T/tau) = exp(-20ns/1us) = exp(-0.02) = 0.9802
        constant C_ALPHA            : real      := 0.9802; -- Matches 1us RC time constant
        variable v_vn               : real      := 0.625;
        variable v_vdac_avg         : real      := 0.0;
        variable v_prev_done        : std_logic := '0';
    begin
        if reset = '1' then
            v_vn             := 0.625;
            analog_voltage_n <= 0.625;
            v_prev_done      := '0';
        elsif rising_edge(clk_tdc) then
            -- Only update on rising edge of duty_period_done
            if duty_period_done = '1' and v_prev_done = '0' then
                v_vdac_avg       := real(duty_count_reg) / real(C_TICKS_PER_PERIOD) * C_DAC_HIGH_V;
                v_vn             := C_ALPHA * v_vn + (1.0 - C_ALPHA) * v_vdac_avg;
                analog_voltage_n <= v_vn;
            end if;
            v_prev_done := duty_period_done;
        end if;
    end process;

    -- ========================================================================
    -- COMPARATOR MODEL - Time-based mode switching for 50MHz reference
    -- ========================================================================
    -- This model serves two distinct purposes:
    -- 
    -- 1. SWEEP MODE (t < 70us): Static comparison for boot sweep detection
    --    - Output reflects instantaneous Vp > Vn comparison
    --    - Required for boot sweep to find crossing duty cycle
    --
    -- 2. TDC MODE (t >= 70us): Generate crossing for TDC measurement
    --    - At ref_clock edge: output starts LOW
    --    - At calculated crossing time: output transitions HIGH
    --    - Crossing time = 8ns + GAIN * (Vp - Vn) for 50MHz (20ns period)
    --    - TDC measures this transition time to generate sample
    p_comparator_model : process
        constant C_SWEEP_END_TIME : time      := 70 us; -- Sweep ends around this time
        variable v_verr           : real      := 0.0; -- Voltage error (Vp - Vn)
        variable v_cross_ns       : real      := 250.0; -- Crossing time in ns
        variable v_pulse_count    : integer   := 0;
        variable v_in_sweep       : boolean   := true; -- True during sweep phase
        variable v_final          : std_logic := '0'; -- Final state for this period
    begin
        -- Initial state before reset
        pad_p <= '0';
        pad_n <= '1';

        wait until reset = '0';

        -- Wait for first ref_clock edge
        wait until rising_edge(ref_clock);

        loop
            -- Sample voltage error at start of period
            v_verr        := analog_voltage_p - analog_voltage_n;
            v_pulse_count := v_pulse_count + 1;

            -- TIME-BASED mode selection (not voltage-based!)
            -- Sweep runs for first ~70us, then closed-loop takes over
            v_in_sweep := now < C_SWEEP_END_TIME;

            if v_in_sweep then
                -- SWEEP MODE: Static output based on voltage comparison
                -- Used during sweep to find crossing duty cycle
                if v_verr > 0.0 then
                    pad_p <= '1';
                    pad_n <= '0';
                else
                    pad_p <= '0';
                    pad_n <= '1';
                end if;

                -- Wait for next ref_clock (no transition needed in sweep mode)
                wait until rising_edge(ref_clock);
            else
                -- ========================================================================
                -- CLOSED LOOP MODE: Delta-sigma feedback with TDC timing info
                -- ========================================================================
                -- Determine final state based on voltage comparison (NOT dac_out_bit!)
                -- This is the delta-sigma comparator decision: Vp > Vn?
                if v_verr > 0.0 then
                    v_final := '1';     -- Vp > Vn: comparator output should be HIGH
                else
                    v_final := '0';     -- Vp <= Vn: comparator output should be LOW
                end if;

                -- For 50MHz (20ns period):
                -- Base offset: 8ns (midpoint of measurement window)
                -- Gain: 3ns/V gives +/-4ns range for +/-1.25V full scale
                -- Result range: 2ns to 18ns (within 20ns period)
                v_cross_ns := 8.0 + (3.0 * v_verr);

                -- Clamp to valid range (must be within reference period)
                if v_cross_ns < 2.0 then
                    v_cross_ns := 2.0;
                elsif v_cross_ns > 18.0 then
                    v_cross_ns := 18.0;
                end if;

                -- Pulse Generation:
                -- 1. Start with opposite state (setup for transition)
                --    Immediate at rising edge (0ns)
                pad_p <= not v_final;
                pad_n <= v_final;

                -- 2. Scheduled transition to final state (measurement edge)
                --    Happens at v_cross_ns after period start
                --    TDC captures this transition BEFORE DAC updates
                pad_p <= transport v_final after v_cross_ns * 1 ns;
                pad_n <= transport not v_final after v_cross_ns * 1 ns;

                -- Wait for next period (Rising Edge)
                wait until rising_edge(ref_clock);
            end if;
        end loop;
    end process;

    -- ========================================================================
    -- RC ADC COMPARATOR MODEL - Simple analog comparison for RC delta-sigma
    -- ========================================================================
    -- For RC ADC, we need a simpler model:
    -- 1. Comparator just compares Vp (input) vs Vn (filtered DAC output)
    -- 2. RC filter models the external capacitor integration of DAC output
    -- 3. No timing-encoded transitions - just instantaneous comparison
    -- ========================================================================

    p_rc_comparator_model : process(clk_sys, reset)
        -- RC filter for DAC feedback modeling at clk_sys rate
        -- Models external RC integrator: DAC_OUT -> R -> C -> ANALOG_IN_N
        constant C_DAC_HIGH_V   : real    := 1.25; -- DAC high voltage (effective Vref)
        constant C_ALPHA        : real    := 0.95; -- RC filter coefficient (~2us time constant at 100MHz)
        variable v_dac_filtered : real    := 0.0; -- Start at 0V to allow proper settling
        variable v_dac_voltage  : real    := 0.0;
        variable v_cycle_count  : integer := 0;
    begin
        if reset = '1' then
            rc_comparator_out <= '0';
            v_dac_filtered    := 0.0;   -- Start at 0V
            v_cycle_count     := 0;
        elsif rising_edge(clk_sys) then
            v_cycle_count := v_cycle_count + 1;

            -- Update DAC filtered voltage
            if dac_out_bit = '1' then
                v_dac_voltage := C_DAC_HIGH_V;
            else
                v_dac_voltage := 0.0;
            end if;

            -- First-order IIR low-pass filter (models RC integration)
            v_dac_filtered := C_ALPHA * v_dac_filtered + (1.0 - C_ALPHA) * v_dac_voltage;

            -- Comparator: Compare input voltage vs filtered DAC output
            if analog_voltage_p > v_dac_filtered then
                rc_comparator_out <= '1';
            else
                rc_comparator_out <= '0';
            end if;
        end if;
    end process;

    -- ========================================================================
    -- Test Runner
    -- ========================================================================
    p_main : process
        -- Convert voltage (0.0-1.0 normalized) to expected Q15 value
        -- V_REF = 1.25V (measured effective reference voltage)
        -- Q15 maps linearly: 0mV -> -32768, 625mV -> 0, 1250mV -> +32767
        -- So: Q15 = (V_normalized - 0.5) * 65536
        function voltage_to_q15(v_normalized : real) return integer is
            variable v_q15 : integer;
        begin
            -- v_normalized is 0.0 to 1.0, mapping to 0mV to 1250mV
            -- Center is 0.5 (625mV) which maps to Q15 = 0
            v_q15 := integer((v_normalized - 0.5) * 65536.0);
            -- Saturate to Q15 range
            if v_q15 > 32767 then
                return 32767;
            elsif v_q15 < -32768 then
                return -32768;
            else
                return v_q15;
            end if;
        end function;

        -- Convert Q15 signed value to millivolts (for reporting only)
        -- V_REF = 1.25V, so center = 625mV, half-scale = 625mV
        -- Formula: mV = (q_value * 625) / 32768 + 625
        -- Q15: -32768 -> 0mV, 0 -> 625mV, +32767 -> 1250mV
        function q_to_mv(q_value : integer) return integer is
            variable v_scaled : integer;
        begin
            -- Scale: multiply by 625, divide by 32768 (2^15)
            v_scaled := (q_value * 625) / 32768 + 625;
            -- Saturate to 0..1250 mV range
            if v_scaled < 0 then
                return 0;
            elsif v_scaled > 1250 then
                return 1250;
            else
                return v_scaled;
            end if;
        end function;

        -- Helper: wait for N sample_valid pulses (deterministic) with timeout and progress monitoring
        procedure wait_for_samples(signal   clk     : std_logic;
                                   signal   vld     : std_logic;
                                   constant N       : natural;
                                   constant timeout : time) is
            variable v_cnt              : unsigned(15 downto 0) := (others => '0');
            variable v_start_time       : time;
            variable v_last_sample_time : time;
            variable v_progress_timer   : time;
        begin
            v_start_time       := now;
            v_last_sample_time := now;
            v_progress_timer   := now;

            while to_integer(v_cnt) < N loop
                wait until rising_edge(clk);

                if vld = '1' then
                    v_cnt              := v_cnt + 1;
                    v_last_sample_time := now;
                    -- Only report progress every 10 samples to reduce output
                    if (to_integer(v_cnt) mod 10) = 0 or to_integer(v_cnt) = N then
                        info("Progress: Collected sample " & integer'image(to_integer(v_cnt)) & " of " & integer'image(N) & " at " & time'image(now));
                    end if;
                end if;

                -- Progress timeout - report if no samples for too long (reduce frequency)
                if now - v_progress_timer > 500 us then
                    info("PROGRESS CHECK: " & integer'image(to_integer(v_cnt)) & " samples collected so far at " & time'image(now) & " (last sample at " & time'image(v_last_sample_time) & ", gap=" & time'image(now - v_last_sample_time) & ")");
                    v_progress_timer := now;
                end if;

                -- Global timeout check
                if now - v_start_time > timeout then
                    error("GLOBAL TIMEOUT waiting for samples! Only got " & integer'image(to_integer(v_cnt)) & " of " & integer'image(N) & " - Last sample at: " & time'image(v_last_sample_time));
                    exit;
                end if;
            end loop;

            info("Sample collection completed: " & integer'image(to_integer(v_cnt)) & " samples in " & time'image(now - v_start_time));
        end procedure;

        -- Helper: Collect samples and verify they are not stuck at zero
        procedure collect_and_verify_samples(signal   clk       : std_logic;
                                             signal   vld       : std_logic;
                                             constant N         : natural;
                                             constant timeout   : time;
                                             constant test_name : string) is
            variable v_mean_mv      : integer;
            variable v_variation_mv : integer;
            variable v_expected_mv  : integer;
            variable v_error_mv     : integer;
            variable v_min_mv       : integer;
            variable v_max_mv       : integer;
            variable v_avg_q        : integer;
            -- Q-format comparison variables
            variable v_expected_q   : integer; -- Expected Q15 value
            variable v_tolerance_q  : integer; -- Tolerance in Q15 units
            variable v_error_q      : integer; -- Error in Q15 units
        begin
            -- Wait for samples to be collected
            wait_for_samples(clk, vld, N, timeout);

            -- Wait for monitoring process to update signals
            wait for C_CLK_SYS_PERIOD * 10;

            -- Check if output is stuck at zero (CRITICAL: This detects broken ADC)
            check(sample_min_value /= 0 or sample_max_value /= 0,
                  "OUTPUT STUCK AT ZERO in " & test_name & ": " & "All " & integer'image(sample_count_sig) & " samples are zero! " & "ADC is not responding to input voltage. " & "Likely causes: " & "1) TDC not generating bitstream " & "2) CIC input stuck " & "3) Servo or mV conversion broken");

            -- Check if output is stuck at constant value (only fail for AC signals)
            -- For DC inputs (GC_TB_SIGNAL_TYPE=1), constant output is expected and correct
            if sample_min_value = sample_max_value and sample_count_sig > 10 and GC_TB_SIGNAL_TYPE /= 1 then
                check(false,
                      "OUTPUT STUCK AT CONSTANT in " & test_name & ": " & "All " & integer'image(sample_count_sig) & " samples equal " & integer'image(sample_min_value) & ". " & "No dynamic range detected for AC signal! Check if: " & "1) Loop is saturated or stuck " & "2) CIC decimation removing all signal variations");
            elsif GC_TB_SIGNAL_TYPE = 1 then
                -- DC INPUT TEST: Verify voltage accuracy in Q15 format
                v_avg_q := sample_sum_value / sample_count_sig; -- Average in Q15

                -- Calculate expected Q15 value from DC level
                -- voltage_to_q15 maps: 0.0 -> -32768, 0.5 -> 0, 1.0 -> +32767
                v_expected_q := voltage_to_q15(GC_TB_DC_LEVEL);

                -- Define tolerance in Q15 units
                -- TDC ADC: +/-10mV corresponds to +/-503 Q15 units (10 * 32768 / 650)
                -- RC ADC: +/-25mV corresponds to +/-1260 Q15 units (25 * 32768 / 650)
                if GC_ADC_TYPE = "rc" then
                    v_tolerance_q := 1260; -- +/-25mV equivalent in Q15
                else
                    v_tolerance_q := 503; -- +/-10mV equivalent in Q15
                end if;
                v_error_q := abs (v_avg_q - v_expected_q);

                -- Convert to mV for reporting only (not for comparison)
                v_min_mv       := q_to_mv(sample_min_value);
                v_max_mv       := q_to_mv(sample_max_value);
                v_mean_mv      := q_to_mv(v_avg_q);
                v_expected_mv  := integer(GC_TB_DC_LEVEL * 1250.0);
                v_variation_mv := v_max_mv - v_min_mv;
                v_error_mv     := abs (v_mean_mv - v_expected_mv);

                -- Report both Q-format and mV values
                info("DC INPUT TEST (Q15): Raw Q15 range " & integer'image(sample_min_value) & " to " & integer'image(sample_max_value) & " (avg=" & integer'image(v_avg_q) & " from " & integer'image(sample_count_sig) & " samples)");
                info("DC INPUT TEST (mV):  Converted range " & integer'image(v_min_mv) & "-" & integer'image(v_max_mv) & "mV (variation=" & integer'image(v_variation_mv) & "mV, avg=" & integer'image(v_mean_mv) & "mV)");
                info("DC ACCURACY (Q15): Expected=" & integer'image(v_expected_q) & ", Measured=" & integer'image(v_avg_q) & ", Error=" & integer'image(v_error_q) & " (tolerance=+/-" & integer'image(v_tolerance_q) & ")");
                info("DC ACCURACY (mV):  Expected=" & integer'image(v_expected_mv) & "mV, Measured=" & integer'image(v_mean_mv) & "mV, Error=" & integer'image(v_error_mv) & "mV");

                -- Check voltage accuracy in Q15 format
                check(v_error_q <= v_tolerance_q,
                      "DC VOLTAGE ERROR EXCEEDS TOLERANCE in " & test_name & ": " & "Expected Q15=" & integer'image(v_expected_q) & " (+/-" & integer'image(v_tolerance_q) & "), " & "Measured Q15=" & integer'image(v_avg_q) & ", " & "Error = " & integer'image(v_error_q) & ". " & "Input voltage: " & integer'image(integer(GC_TB_DC_LEVEL * 1250.0)) & "mV.");

                info("DC VOLTAGE ACCURACY CHECK PASSED: Error Q15=" & integer'image(v_error_q) & " within +/-" & integer'image(v_tolerance_q) & " tolerance");
            else
                -- For AC signals (sine, square, ramp), just verify dynamic range exists
                -- The ADC outputs absolute voltage (0-1200mV), not differential amplitude
                -- So for a 0.25 amplitude sine at 0.5 DC offset (300mV swing centered at 600mV),
                -- the output range will be close to full scale as the loop tracks the input
                v_min_mv       := q_to_mv(sample_min_value);
                v_max_mv       := q_to_mv(sample_max_value);
                v_variation_mv := v_max_mv - v_min_mv; -- Peak-to-peak in mV

                info("AC INPUT TEST (Q15): Raw Q15 range " & integer'image(sample_min_value) & " to " & integer'image(sample_max_value));
                info("AC INPUT TEST (mV):  Peak-to-peak range = " & integer'image(v_variation_mv) & " mV (" & integer'image(v_min_mv) & "-" & integer'image(v_max_mv) & "mV)");

                -- Just verify we have reasonable dynamic range (>100mV) to confirm loop is tracking
                check(v_variation_mv > 100,
                      "AC OUTPUT HAS NO DYNAMIC RANGE in " & test_name & ": " & "Only " & integer'image(v_variation_mv) & "mV p-p detected " & "(AMPLITUDE=" & real'image(GC_TB_AMPLITUDE) & ", FREQUENCY=" & real'image(GC_TB_FREQUENCY_HZ) & "Hz). " & "Delta-Sigma loop may be stuck!");

                info("AC VOLTAGE TRACKING CHECK PASSED: Measured " & integer'image(v_variation_mv) & "mV p-p dynamic range");
            end if;

            info("OUTPUT RANGE CHECK PASSED for " & test_name & ": Q15 min=" & integer'image(sample_min_value) & ", max=" & integer'image(sample_max_value) & ", count=" & integer'image(sample_count_sig));
        end procedure;

    begin
        test_runner_setup(runner, runner_cfg);

        while test_suite loop
            if run("basic_test") then
                info("==========================================================");
                info("Running TDC ADC basic test with external analog input");
                info("Signal type: " & integer'image(GC_TB_SIGNAL_TYPE));
                info("DC level: " & real'image(GC_TB_DC_LEVEL));
                info("Amplitude: " & real'image(GC_TB_AMPLITUDE));
                info("Frequency: " & real'image(GC_TB_FREQUENCY_HZ) & " Hz");
                info("==========================================================");

                -- DYNAMIC READY DETECTION: Wait for first sample_valid pulse
                -- This indicates calibration is complete and system is producing valid output
                info("Waiting for system ready (first sample_valid)...");
                wait until rising_edge(clk_sys) and sample_valid = '1' for 500 us;
                if sample_valid /= '1' then
                    error("Timeout waiting for first sample_valid - calibration may have failed!");
                end if;
                info("System ready detected at " & time'image(now));

                -- Collect samples for accuracy measurement
                -- TDC @ 2MHz -> Decimation /64 -> ~31.25kHz (~32us period)
                -- RC @ 100MHz -> Decimation /64 -> ~1.5625MHz (~640ns period)
                -- RC ADC needs ~120 samples for FIR filter priming (31+63 taps + margin)
                -- After priming, need additional samples for measurement
                if GC_TB_SIGNAL_TYPE = 1 then
                    -- DC test
                    if GC_ADC_TYPE = "rc" then
                        -- RC ADC: 125 samples (120 settling + 5 measurement), ~80us at 1.5MHz
                        info("Collecting 125 output samples for RC ADC DC accuracy test (120 settling + 5 measurement)...");
                        collect_and_verify_samples(clk_sys, sample_valid, 125, 200 us, "basic_test");
                    else
                        -- TDC ADC: 75 samples (70 filter priming + 5 measurement), 2.5ms timeout
                        -- Filter priming count is 70 samples before combined CIC/EQ/LP+TDC output is stable
                        -- 75 samples @ 32us each = 2.4ms - use 2.5ms timeout
                        info("Collecting 75 output samples for TDC ADC DC accuracy test (70 settling + 5 measurement)...");
                        collect_and_verify_samples(clk_sys, sample_valid, 75, 2500 us, "basic_test");
                    end if;
                else
                    -- AC test (sine/square/ramp)
                    if GC_ADC_TYPE = "rc" then
                        -- RC ADC: 220 samples (120 settling + 100 measurement)
                        info("Collecting 220 output samples for RC ADC AC test (120 settling + 100 measurement)...");
                        collect_and_verify_samples(clk_sys, sample_valid, 220, 500 us, "basic_test");
                    else
                        -- TDC ADC: 100 samples, 25ms timeout
                        info("Collecting 100 output samples for TDC ADC AC test (includes filter priming)...");
                        collect_and_verify_samples(clk_sys, sample_valid, 100, 25 ms, "basic_test");
                    end if;
                end if;

                info("==========================================================");
                info("Basic test completed successfully");
                info("==========================================================");

            elsif run("digital_self_test") then
                info("==========================================================");
                info("Running TDC ADC DIGITAL SELF-TEST mode (internal digital test signal)");
                info("Note: DUT configured with GC_SELF_TEST=false");
                info("This tests external analog path with time-domain modulation");
                info("In hardware with GC_SELF_TEST=true, both Stop and TDL edge");
                info("are generated internally as DIGITAL pulses for deterministic timing");
                info("==========================================================");

                -- Wait for reset + settle (ADC uses default configuration)
                wait for C_CLK_SYS_PERIOD * 100;

                -- Wait for samples - should work with external analog stimulus
                -- when GC_SELF_TEST=true in hardware, uses internal digital test signals
                -- Timeout calculation: TDC @ 2MHz -> CIC /64 -> ~31.25kHz (32us period)
                -- Need ~63 (FIR fill) + 20 samples = 83 samples x 32us = 2656us = 3ms
                info("Waiting for 20 output samples (digital self-test configuration)...");
                collect_and_verify_samples(clk_sys, sample_valid, 20, 5 ms, "digital_self_test");

                info("==========================================================");
                info("Digital self-test completed - system produces stable output");
                info("Coarse timestamp fix verified in digital self-test mode!");
                info("==========================================================");

            elsif run("tdc_characterization") then
                info("==========================================================");
                info("TDC 2D CHARACTERIZATION TEST - Fast DAC Duty Sweep");
                info("Input Voltage: " & integer'image(integer(GC_TB_DC_LEVEL * 1250.0)) & "mV");
                info("Sweeping DAC duty: 40%, 50%, 60% (3 points around midpoint)");
                info("Goal: Find if ANY region has unsaturated TDC output");
                info("==========================================================");

                -- Wait for reset + settle
                wait for C_CLK_SYS_PERIOD * 100;

                -- Sweep DAC duty from 40% to 60% in 10% increments (3 points)
                -- For each duty, collect TDC statistics until 2000 samples
                for duty_pct in 4 to 6 loop -- 40%, 50%, 60% only
                    -- Pulse testpoint_reset to clear TDC monitor accumulators
                    testpoint_reset <= '1';
                    wait for 1 us;
                    testpoint_reset <= '0';
                    wait for 1 us;

                    info("======================================================");
                    info("Test Point: Vin=" & integer'image(integer(GC_TB_DC_LEVEL * 1250.0)) & "mV, DAC=" & integer'image(duty_pct * 10) & "%");
                    info("Expected Vdac_avg ~= " & integer'image(duty_pct * 125) & "mV");
                    info("Expected differential ~= " & integer'image(integer(GC_TB_DC_LEVEL * 1250.0) - duty_pct * 125) & "mV");

                    -- Generate PWM at ref_clock rate (2 MHz = 500ns period)
                    -- duty_pct=4..6 -> PWM with 40%, 50%, 60% duty cycle
                    -- Wait until tdc_char_done (2000 samples) instead of fixed 5ms

                    -- Reset TDC monitor stats via testpoint_reset pulse
                    -- This also resets tdc_char_done in p_tdc_monitor
                    testpoint_reset <= '1';
                    wait for 100 ns;
                    testpoint_reset <= '0';
                    wait for 100 ns;

                    -- PWM: Toggle at ref_clock rate with specified duty cycle
                    -- ref period = 500ns, so high time = duty_pct * 50ns
                    -- Loop until 2000 TDC samples collected (tdc_char_done = true)
                    while not tdc_char_done loop
                        open_loop_dac <= '1';
                        wait for (duty_pct * 50) * 1 ns;
                        open_loop_dac <= '0';
                        wait for ((10 - duty_pct) * 50) * 1 ns;
                    end loop;

                    info("Completed measurement at " & integer'image(duty_pct * 10) & "% duty");
                end loop;

                info("==========================================================");
                info("2D Characterization completed - 3 DAC duties tested (40-60%)");
                info("Analyze TDC_LOG output to find usable operating regions");
                info("==========================================================");

            elsif run("pi_step_response") then
                -- ============================================================
                -- PI STEP RESPONSE TEST - Closed-loop tuning
                -- ============================================================
                -- This test is for tuning PI gains with GC_OPEN_LOOP=false
                -- 1. Start at mid-scale (GC_TB_DC_LEVEL), let loop settle
                -- 2. Step input to GC_TB_DC_LEVEL + 0.1 (130mV step)
                -- 3. Measure settling time, overshoot, oscillation
                -- ============================================================
                info("==========================================================");
                info("PI STEP RESPONSE TEST - Closed-Loop Tuning");
                info("Initial DC level: " & real'image(GC_TB_DC_LEVEL));
                info("NOTE: Must run with GC_OPEN_LOOP=false for closed-loop!");
                info("==========================================================");

                -- Wait for reset + calibration + initial settling
                info("Phase 1: Waiting for boot + calibration (~200us)...");
                wait for 200 us;

                -- Let loop settle at initial operating point
                info("Phase 2: Initial settling at " & real'image(GC_TB_DC_LEVEL) & " for 500us...");
                wait for 500 us;

                info("Phase 3: Collecting samples to measure settling behavior...");

                -- Reset sample statistics
                testpoint_reset <= '1';
                wait for 100 ns;
                testpoint_reset <= '0';

                -- Collect samples for 1ms and observe statistics
                collect_and_verify_samples(clk_sys, sample_valid, 100, 5 ms, "pi_step_response");

                info("==========================================================");
                info("PI Step Response test completed");
                info("Check RC_AVG and PI_LOOP logs for settling behavior");
                info("==========================================================");

            end if;
        end loop;

        wait for C_CLK_SYS_PERIOD * 10;
        sim_finished <= true;
        test_runner_cleanup(runner);
        wait;
    end process;

    -- ========================================================================
    -- Sample Monitor
    -- ========================================================================
    -- SETTLING SAMPLE THRESHOLD: Discard early transient samples from DC statistics
    -- The delta-sigma loop needs time to settle after boot. Early samples during
    -- SWEEP/DITHER/early closed-loop will have large errors and should not be
    -- included in DC accuracy calculations. Only samples AFTER this threshold
    -- are used for min/max/avg statistics.
    -- 
    -- With FIR lowpass filter (63 taps), need 63+ samples to fill delay line.
    -- Add extra margin for CIC/equalizer/PI loop settling.
    -- RC ADC needs more settling due to 31-tap EQ + 63-tap LP = 94 taps total

    p_monitor : process(clk_sys)
        -- RC ADC needs more settling due to FIR filter delay lines (31 + 63 = 94 taps)
        -- TDC ADC has filter priming count of 70 samples before combined output is stable
        -- Add margin: RC needs ~120 samples, TDC needs ~70
        constant C_SETTLE_SAMPLES_TDC : integer := 70; -- Match C_FILTER_PRIME_COUNT in tdc_adc_top
        constant C_SETTLE_SAMPLES_RC  : integer := 120; -- 94 taps + margin
        variable v_settle_limit       : integer;
        variable v_sample_count       : integer := 0; -- Total samples seen (including settling)
        variable v_stats_count        : integer := 0; -- Samples used for statistics (after settling)
        variable v_min_value          : integer := integer'high;
        variable v_max_value          : integer := integer'low;
        variable v_sum                : integer := 0;
        variable v_sample_value       : integer;
    begin
        if rising_edge(clk_sys) then
            -- Select settling limit based on ADC type
            if GC_ADC_TYPE = "rc" then
                v_settle_limit := C_SETTLE_SAMPLES_RC;
            else
                v_settle_limit := C_SETTLE_SAMPLES_TDC;
            end if;

            if reset = '1' then
                v_sample_count   := 0;
                v_stats_count    := 0;
                v_min_value      := integer'high;
                v_max_value      := integer'low;
                v_sum            := 0;
                sample_min_value <= 0;
                sample_max_value <= 0;
                sample_count_sig <= 0;
                sample_sum_value <= 0;
            elsif sample_valid = '1' then
                v_sample_count := v_sample_count + 1;
                v_sample_value := to_integer(signed(sample_data));

                -- Only include samples AFTER settling period in statistics
                if v_sample_count > v_settle_limit then
                    v_stats_count := v_stats_count + 1;
                    v_sum         := v_sum + v_sample_value;

                    -- Track min/max (only settled samples)
                    if v_sample_value < v_min_value then
                        v_min_value := v_sample_value;
                    end if;
                    if v_sample_value > v_max_value then
                        v_max_value := v_sample_value;
                    end if;
                end if;

                -- Update signals for test process to check (only after settling)
                if v_sample_count > v_settle_limit and v_stats_count > 0 then
                    sample_min_value <= v_min_value;
                    sample_max_value <= v_max_value;
                    sample_count_sig <= v_stats_count; -- Report settled sample count
                    sample_sum_value <= v_sum;
                end if;

                -- Reduced debug output for speed - only print first 5 and last sample
                if v_sample_count <= 5 then
                    info("Sample " & integer'image(v_sample_count) & " [SETTLING]: " & integer'image(v_sample_value));
                elsif v_sample_count = v_settle_limit + 1 then
                    info("=== SETTLING COMPLETE (" & integer'image(v_settle_limit) & " samples discarded) ===");
                end if;
            end if;
        end if;
    end process;

    -- ========================================================================
    -- TDC Monitor - Enhanced statistics for 2D characterization
    -- With early termination support: sets tdc_char_done after 2000 samples
    -- Only enabled for characterization tests (GC_OPEN_LOOP=true)
    -- ========================================================================
    g_tdc_monitor : if GC_OPEN_LOOP generate
        p_tdc_monitor : process(clk_tdc)
            variable v_tdc_count          : integer := 0;
            variable v_tdc_sum            : integer := 0;
            variable v_tdc_sum_sq         : integer := 0; -- Sum of squares for stddev
            variable v_tdc_min            : integer := integer'high;
            variable v_tdc_max            : integer := integer'low;
            variable v_tdc_sat_count      : integer := 0; -- Count of saturated samples (+/-128)
            variable v_tdc_value          : integer;
            variable v_mean               : integer;
            variable v_variance           : integer;
            variable v_sat_pct            : integer;
            constant C_CHAR_SAMPLE_TARGET : integer := 2000; -- Early termination threshold
        begin
            if rising_edge(clk_tdc) then
                -- Reset on global reset OR testpoint_reset pulse
                if reset = '1' or testpoint_reset = '1' then
                    v_tdc_count     := 0;
                    v_tdc_sum       := 0;
                    v_tdc_sum_sq    := 0;
                    v_tdc_min       := integer'high;
                    v_tdc_max       := integer'low;
                    v_tdc_sat_count := 0;
                    tdc_char_done   <= false; -- Reset early termination flag
                elsif debug_tdc_valid = '1' and not tdc_char_done then
                    v_tdc_value  := to_integer(debug_tdc_out);
                    v_tdc_count  := v_tdc_count + 1;
                    v_tdc_sum    := v_tdc_sum + v_tdc_value;
                    v_tdc_sum_sq := v_tdc_sum_sq + (v_tdc_value * v_tdc_value);

                    -- Track saturation: TDC saturates when coarse count hits limits
                    -- With 8-bit coarse counter and 8 fractional bits, saturation is:
                    --   Max positive: +(2^7 - 1) x 256 = +32512 codes
                    --   Max negative: -(2^7) x 256 = -32768 codes
                    -- Use conservative threshold of +/-30000 to detect approaching saturation
                    if abs (v_tdc_value) >= 30000 then
                        v_tdc_sat_count := v_tdc_sat_count + 1;
                    end if;

                    if v_tdc_value < v_tdc_min then
                        v_tdc_min := v_tdc_value;
                    end if;
                    if v_tdc_value > v_tdc_max then
                        v_tdc_max := v_tdc_value;
                    end if;

                    -- Log every 2000th sample with full statistics (reduced for speed)
                    if (v_tdc_count mod 2000) = 0 then
                        v_mean     := v_tdc_sum / v_tdc_count;
                        v_variance := (v_tdc_sum_sq / v_tdc_count) - (v_mean * v_mean);
                        v_sat_pct  := (v_tdc_sat_count * 100) / v_tdc_count;

                        info("TDC_STAT: n=" & integer'image(v_tdc_count) & " mean=" & integer'image(v_mean) & " var=" & integer'image(v_variance) & " range=[" & integer'image(v_tdc_min) & "," & integer'image(v_tdc_max) & "]" & " sat=" & integer'image(v_sat_pct) & "%" & " Vin=" & integer'image(integer(analog_voltage_p * 1000.0)) & "mV" & " Vdac=" & integer'image(integer(analog_voltage_n * 1000.0)) & "mV" & " dV=" & integer'image(integer((analog_voltage_p - analog_voltage_n) * 1000.0)) & "mV" & " DAC=" & std_logic'image(open_loop_dac));
                    end if;

                    -- Early termination: signal done after reaching sample target
                    if v_tdc_count >= C_CHAR_SAMPLE_TARGET then
                        tdc_char_done <= true;
                    end if;
                end if;
            end if;
        end process;
    end generate g_tdc_monitor;

    -- ========================================================================
    -- Watchdog Monitor - Reports system status periodically (disabled for speed)
    -- ========================================================================
    p_watchdog : process
        constant C_REPORT_INTERVAL : time := 1 ms; -- Increased from 100us for speed
    begin
        wait until reset = '0';

        loop
            wait for C_REPORT_INTERVAL;

            if not sim_finished then
                info("WATCHDOG at " & time'image(now) & " sample_data=" & integer'image(to_integer(signed(sample_data))));
            else
                exit;
            end if;
        end loop;
        wait;
    end process;

end architecture behavioral;
