-- ************************************************************************
-- Simplified Delta-Sigma ADC Top Level for AXE5000
-- Minimal integration with NIOS-V using Avalon-MM interface
-- ************************************************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Note: library work is implicit, no need to declare
use work.clk_rst_pkg.all;

entity axe5000_top is
  generic(
    ADC_DECIMATION : positive := 64     -- Configurable OSR/decimation factor
  );
  port(
    -- Clock and Reset
    CLK_25M_C  : in  std_logic;
    CPU_RESETn : in  std_logic;
    -- UART
    UART_TX    : out std_logic;
    UART_RX    : in  std_logic;
    -- DIP Switches
    DIP_SW     : in  std_logic_vector(1 downto 0);
    -- Delta-Sigma ADC (differential LVDS input)
    ANALOG_IN  : in  std_logic;         -- From comparator (differential pair handled at I/O level)
    DAC_OUT    : out std_logic;         -- To integrator/filter

    -- Debug
    TEST_PIN   : out std_logic
  );
end entity;

architecture rtl of axe5000_top is

  signal clk_100m     : std_logic;
  signal reset_n      : std_logic;
  signal system_reset : rst_t;

  -- Clock crossing bridge signals
  signal bridge_clk           : std_logic;
  signal bridge_reset         : std_logic;
  signal bridge_waitrequest   : std_logic;
  signal bridge_readdata      : std_logic_vector(31 downto 0);
  signal bridge_readdatavalid : std_logic;
  signal bridge_writedata     : std_logic_vector(31 downto 0);
  signal bridge_address       : std_logic_vector(15 downto 0);
  signal bridge_write         : std_logic;
  signal bridge_read          : std_logic;

  -- Address decoder signals
  constant NUM_MODULES       : natural := 2; -- ADC + About
  signal   mem_cs            : std_logic_vector(NUM_MODULES - 1 downto 0);
  signal   mem_rd            : std_logic;
  signal   mem_wr            : std_logic;
  signal   mem_addr          : std_logic_vector(11 downto 0); -- 12-bit for 4KB range
  signal   mem_wdata         : std_logic_vector(31 downto 0);
  signal   mem_rdata_array_0 : std_logic_vector(31 downto 0); -- ADC module
  signal   mem_rdata_array_1 : std_logic_vector(31 downto 0); -- About module
  signal   mem_rdvalid       : std_logic_vector(NUM_MODULES - 1 downto 0);

  -- ADC module signals
  signal adc_rdata   : std_logic_vector(31 downto 0);
  signal adc_rdvalid : std_logic;

  -- About module signals  
  signal about_rdata   : std_logic_vector(31 downto 0);
  signal about_rdvalid : std_logic;

  -- NIOS-V system component (generated by Platform Designer)
  component niosv_system is             -- @suppress
    port(
      clk_25m_clk               : in  std_logic;
      dip_sw_export             : in  std_logic_vector(1 downto 0);
      uart_rxd                  : in  std_logic;
      uart_txd                  : out std_logic;
      mm_ccb_0_m0_clk_clk       : in  std_logic;
      mm_ccb_0_m0_reset_reset   : in  std_logic;
      mm_ccb_0_m0_waitrequest   : in  std_logic;
      mm_ccb_0_m0_readdata      : in  std_logic_vector(31 downto 0);
      mm_ccb_0_m0_readdatavalid : in  std_logic;
      mm_ccb_0_m0_burstcount    : out std_logic_vector(0 downto 0);
      mm_ccb_0_m0_writedata     : out std_logic_vector(31 downto 0);
      mm_ccb_0_m0_address       : out std_logic_vector(15 downto 0);
      mm_ccb_0_m0_write         : out std_logic;
      mm_ccb_0_m0_read          : out std_logic;
      mm_ccb_0_m0_byteenable    : out std_logic_vector(3 downto 0);
      mm_ccb_0_m0_debugaccess   : out std_logic;
      reset_n_reset_n           : in  std_logic;
      sysclk_clk                : out std_logic
    );
  end component;

begin

  -- Reset management
  reset_n      <= CPU_RESETn;
  system_reset <= not reset_n;

  -- Debug output
  TEST_PIN <= ANALOG_IN;                -- Simple debug signal

  -- Bridge clock domain uses the 100MHz system clock
  bridge_clk   <= clk_100m;
  bridge_reset <= system_reset;

  -- NIOS-V System with Clock Crossing Bridge
  niosv_inst : niosv_system
    port map(
      clk_25m_clk               => CLK_25M_C,
      dip_sw_export             => DIP_SW,
      uart_rxd                  => UART_RX,
      uart_txd                  => UART_TX,
      mm_ccb_0_m0_clk_clk       => bridge_clk,
      mm_ccb_0_m0_reset_reset   => bridge_reset,
      mm_ccb_0_m0_waitrequest   => bridge_waitrequest,
      mm_ccb_0_m0_readdata      => bridge_readdata,
      mm_ccb_0_m0_readdatavalid => bridge_readdatavalid,
      mm_ccb_0_m0_burstcount    => open, -- Not used for simple peripherals
      mm_ccb_0_m0_writedata     => bridge_writedata,
      mm_ccb_0_m0_address       => bridge_address,
      mm_ccb_0_m0_write         => bridge_write,
      mm_ccb_0_m0_read          => bridge_read,
      mm_ccb_0_m0_byteenable    => open, -- Not used for word-aligned access
      mm_ccb_0_m0_debugaccess   => open,
      reset_n_reset_n           => reset_n,
      sysclk_clk                => clk_100m
    );

  -- Address Decoder: Routes bridge requests to ADC/About modules
  addr_decoder_inst : entity work.addr_decoder
    generic map(
      GC_BRIDGE_ADDR_W => 16,
      GC_MEM_DATA_W    => 32,
      GC_MEM_ADDR_W    => 12,
      GC_NUM_MODULES   => NUM_MODULES
    )
    port map(
      clk               => bridge_clk,
      bridge_rd         => bridge_read,
      bridge_wr         => bridge_write,
      bridge_addr       => bridge_address,
      bridge_wdata      => bridge_writedata,
      bridge_rdata      => bridge_readdata,
      bridge_rdvalid    => bridge_readdatavalid,
      mem_cs            => mem_cs,
      mem_rd            => mem_rd,
      mem_wr            => mem_wr,
      mem_addr          => mem_addr,
      mem_wdata         => mem_wdata,
      mem_rdata_array_0 => mem_rdata_array_0,
      mem_rdata_array_1 => mem_rdata_array_1,
      mem_rdvalid       => mem_rdvalid
    );

  -- Bridge waitrequest (no wait states for simple modules)
  bridge_waitrequest <= '0';

  -- Connect individual module read data to array
  mem_rdata_array_0 <= adc_rdata;       -- ADC module
  mem_rdata_array_1 <= about_rdata;     -- About module
  mem_rdvalid       <= (0 => adc_rdvalid, 1 => about_rdvalid);

  -- ADC Module (placeholder - connect to your rc_adc_top)
  adc_inst : entity work.rc_adc_top
    generic map(
      DECIMATION      => ADC_DECIMATION,
      DATA_WIDTH      => 16,
      ENABLE_MAJORITY => false
    )
    port map(
      clk         => bridge_clk,
      reset       => bridge_reset,
      -- Memory interface
      mem_cs      => mem_cs(0),         -- ADC module index
      mem_rd      => mem_rd,
      mem_wr      => mem_wr,
      mem_addr    => mem_addr,
      mem_wdata   => mem_wdata,
      mem_rdata   => adc_rdata,
      mem_rdvalid => adc_rdvalid,
      -- ADC interface
      analog_in_p => ANALOG_IN,
      analog_in_n => '0',               -- Not used - differential handled at I/O level
      dac_out     => DAC_OUT
    );

  -- About Module: Provides version and build information
  about_inst : entity work.about
    generic map(
      GC_MEM_ADDR_W      => 12,
      GC_MEM_DATA_W      => 32,
      GC_IMAGE_TYPE      => 1,          -- ADC Project Type
      GC_IMAGE_ID        => 16#5000#,   -- AXE5000 ID
      GC_REV_MAJOR       => 1,          -- Major version
      GC_REV_MINOR       => 0,          -- Minor version  
      GC_REV_PATCH       => 0,          -- Patch version
      GC_REV_BUILDNUMBER => 1,          -- Build number
      GC_GIT_HASH_MSB    => 0,          -- Git hash upper
      GC_GIT_HASH_LSB    => 0,          -- Git hash lower
      GC_GIT_DIRTY       => 0,          -- Git clean
      GC_YYMMDD          => 16#250911#, -- Build date (2025-09-11)
      GC_HHMMSS          => 16#120000#  -- Build time (12:00:00)
    )
    port map(
      clk         => bridge_clk,
      mem_cs      => mem_cs(1),         -- About module index
      mem_rd      => mem_rd,
      mem_addr    => mem_addr,
      mem_rdata   => about_rdata,
      mem_rdvalid => about_rdvalid
    );

end architecture rtl;
